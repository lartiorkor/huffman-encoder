	----------------------------------------------------------------------------------
	-- Company: 
	-- Engineer: 
	-- 
	-- Create Date:    18:36:22 11/29/2021 
	-- Design Name: 
	-- Module Name:    adder - Behavioral 
	-- Project Name: 
	-- Target Devices: 
	-- Tool versions: 
	-- Description: 
	--
	-- Dependencies: 
	--
	-- Revision: 
	-- Revision 0.01 - File Created
	-- Additional Comments: 
	--
	----------------------------------------------------------------------------------
	library IEEE;
	use IEEE.STD_LOGIC_1164.ALL;
	use IEEE.STD_LOGIC_UNSIGNED.ALL;

	-- Uncomment the following library declaration if using
	-- arithmetic functions with Signed or Unsigned values
	use IEEE.NUMERIC_STD.ALL;

	-- Uncomment the following library declaration if instantiating
	-- any Xilinx primitives in this code.
	--library UNISIM;
	--use UNISIM.VComponents.all;

	entity adder is 
	
	Port( 
	data_in_1 : in  std_logic_vector(3 downto 0);
	data_in_2 : in  std_logic_vector(3 downto 0);
	data_out  : out std_logic_vector(3 downto 0)
	);
	
	end adder;

	architecture Behavioral of adder is
	
	begin
	
	data_out <= data_in_1 + data_in_2;


	end Behavioral;

